module f_function (

		output wire [1023:0] v_out,
		input wire clk,
		input [1023:0] v,
		input [1023:0]chunk
	);	
	
	
	wire [64*16-1:0] v_con [0:12*8];

	
	localparam [0:4*8*4-1] v_index = {
  4'd0, 4'd4, 4'd8, 4'd12,
  4'd1, 4'd5, 4'd9, 4'd13,
  4'd2, 4'd6, 4'd10, 4'd14,
  4'd3, 4'd7, 4'd11, 4'd15,

  4'd0, 4'd5, 4'd10, 4'd15,
  4'd1, 4'd6, 4'd11, 4'd12,
  4'd2, 4'd7, 4'd8, 4'd13,
  4'd3, 4'd4, 4'd9, 4'd14
};


	localparam [0:4*16*12-1] SIGMA = {
  4'd0, 4'd1, 4'd2, 4'd3, 4'd4, 4'd5, 4'd6, 4'd7, 4'd8, 4'd9, 4'd10, 4'd11, 4'd12, 4'd13, 4'd14, 4'd15,
  4'd14, 4'd10, 4'd4, 4'd8, 4'd9, 4'd15, 4'd13, 4'd6, 4'd1, 4'd12, 4'd0, 4'd2, 4'd11, 4'd7, 4'd5, 4'd3,
  4'd11, 4'd8, 4'd12, 4'd0, 4'd5, 4'd2, 4'd15, 4'd13, 4'd10, 4'd14, 4'd3, 4'd6, 4'd7, 4'd1, 4'd9, 4'd4,
  4'd7, 4'd9, 4'd3, 4'd1, 4'd13, 4'd12, 4'd11, 4'd14, 4'd2, 4'd6, 4'd5, 4'd10, 4'd4, 4'd0, 4'd15, 4'd8,
  4'd9, 4'd0, 4'd5, 4'd7, 4'd2, 4'd4, 4'd10, 4'd15, 4'd14, 4'd1, 4'd11, 4'd12, 4'd6, 4'd8, 4'd3, 4'd13,
  4'd2, 4'd12, 4'd6, 4'd10, 4'd0, 4'd11, 4'd8, 4'd3, 4'd4, 4'd13, 4'd7, 4'd5, 4'd15, 4'd14, 4'd1, 4'd9,
  4'd12, 4'd5, 4'd1, 4'd15, 4'd14, 4'd13, 4'd4, 4'd10, 4'd0, 4'd7, 4'd6, 4'd3, 4'd9, 4'd2, 4'd8, 4'd11,
  4'd13, 4'd11, 4'd7, 4'd14, 4'd12, 4'd1, 4'd3, 4'd9, 4'd5, 4'd0, 4'd15, 4'd4, 4'd8, 4'd6, 4'd2, 4'd10,
  4'd6, 4'd15, 4'd14, 4'd9, 4'd11, 4'd3, 4'd0, 4'd8, 4'd12, 4'd2, 4'd13, 4'd7, 4'd1, 4'd4, 4'd10, 4'd5,
  4'd10, 4'd2, 4'd8, 4'd4, 4'd7, 4'd6, 4'd1, 4'd5, 4'd15, 4'd11, 4'd9, 4'd14, 4'd3, 4'd12, 4'd13, 4'd0,
  4'd0, 4'd1, 4'd2, 4'd3, 4'd4, 4'd5, 4'd6, 4'd7, 4'd8, 4'd9, 4'd10, 4'd11, 4'd12, 4'd13, 4'd14, 4'd15,
  4'd14, 4'd10, 4'd4, 4'd8, 4'd9, 4'd15, 4'd13, 4'd6, 4'd1, 4'd12, 4'd0, 4'd2, 4'd11, 4'd7, 4'd5, 4'd3
};


	mix mix_r0_0(.clk(clk), .v(v), .a(4'd0), .b(4'd4), .c(4'd8), .d(4'd12), .x(chunk[0*64 +: 64]), .y(chunk[1*64 +: 64]), .v_out(v_con[1]));
	
	generate
	  genvar i;
	  for(i = 1; i < 12*8; i = i + 1)
	  begin: generate_mix_rounds
		 mix mix_rround_i(
			.clk(clk),
			.v(v_con[i]),
			.a(v_index[ ((i*16) + 0)%128+:4 ]),
			.b(v_index[ ((i*16) + 4)%128+:4 ]),
			.c(v_index[ ((i*16) + 8)%128+:4 ]),
			.d(v_index[ ((i*16) + 12)%128+:4 ]),
			.x(chunk[ SIGMA[ i*8 +: 4 ]*64 +: 64]),
			.y(chunk[ SIGMA[ i*8+4 +: 4 ]*64 +: 64]),
			.v_out(v_con[i+1])
		 );
	  end
	endgenerate
	assign v_out = v_con[96];

endmodule